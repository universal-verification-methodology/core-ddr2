/**
 * Icarus Verilog testbench for ddr2_server_controller.
 * Currently exercises the same scenarios as tb_ddr2_controller, but instantiates
 * the server-style top cell (`ddr2_server_controller`) instead of the plain
 * `ddr2_controller`. This keeps the test logic identical while allowing the
 * server wrapper to evolve independently (e.g. wider data paths, multi-rank).
 */
`timescale 1ns/1ps

/* verilator lint_off UNUSEDSIGNAL */
module tb_ddr2_server_controller;

    reg         CLK;
    reg         RESET;
    reg         INITDDR;
    reg  [2:0]  CMD;
    reg  [1:0]  SZ;
    reg  [24:0] ADDR;
    reg         cmd_put;
    // 64-bit host data bus for the server-style top (4×16-bit slices).
    reg  [63:0] DIN;
    reg         put_dataFIFO;
    reg         FETCHING;
    // Optional low-power controls mirrored from the core controller. These are
    // held low for the legacy scenarios and driven only in the dedicated
    // power-management tests.
    reg         SELFREF_REQ;
    reg         SELFREF_EXIT;
    reg         PWRDOWN_REQ;
    reg         PWRDOWN_EXIT;
    // Optional runtime DLL controls for the server top; currently forwarded
    // directly to the underlying core controller slice 0.
    reg         DLL_REQ;
    reg         DLL_MODE;
    wire [63:0] DOUT;
    wire [24:0] RADDR;
    wire [6:0]  FILLCOUNT;
    wire        READY;
    wire        VALIDOUT;
    wire        NOTFULL;
    // Two-rank CS# vector on the DDR2 bus (active low).
    wire [1:0]  C0_CSBAR_PAD;
    wire        C0_RASBAR_PAD;
    wire        C0_CASBAR_PAD;
    wire        C0_WEBAR_PAD;
    wire [1:0]  C0_BA_PAD;
    wire [12:0] C0_A_PAD;
    wire [1:0]  C0_DM_PAD;
    wire        C0_ODT_PAD;
    wire        C0_CK_PAD;
    wire        C0_CKBAR_PAD;
    wire        C0_CKE_PAD;
    wire [15:0] C0_DQ_PAD;
    wire [1:0]  C0_DQS_PAD;
    wire [1:0]  C0_DQSBAR_PAD;

    // Internal variables for checking.
    integer cycle;
    integer i;
    integer csv_fd;
`ifdef NEGATIVE_TESTS
    // Flag used to distinguish intentional illegal commands in NEGATIVE_TESTS
    // from accidental ones during the main positive test phases.
    reg neg_expect_illegal_cmd;
`endif

    // Simple functional coverage counters (per-command and per-SZ).
    integer cov_scw, cov_scr, cov_blw, cov_blr;
    integer cov_sz0, cov_sz1, cov_sz2, cov_sz3;

    // ------------------------------------------------------------------------
    // Data pattern and simple scoreboard for read-back verification.
    // ------------------------------------------------------------------------

    // Deterministic data pattern as a function of address.
    function [15:0] pattern_for_addr;
        input [24:0] addr;
        begin
            pattern_for_addr = {addr[7:0], addr[15:8]} ^ 16'hA5A5;
        end
    endfunction

    // Very simple scoreboard using parallel arrays.
    integer sb_idx;
    integer sb_size;
    reg [24:0] sb_addr [0:2047];
    // Expected 64-bit word per address (4× identical 16-bit lanes).
    reg [63:0] sb_data [0:2047];

    task automatic sb_reset;
        begin
            sb_size = 0;
        end
    endtask

    task automatic sb_write;
        input [24:0] addr;
        input [63:0] data;
        reg          updated;
        begin
            // Overwrite if address already present; otherwise append a new
            // entry. Avoids use of "disable task" so that static analysis
            // tools like Verilator can lint this code.
            updated = 1'b0;
            for (sb_idx = 0; sb_idx < sb_size; sb_idx = sb_idx + 1) begin
                if (sb_addr[sb_idx] == addr) begin
                    sb_data[sb_idx] = data;
                    updated = 1'b1;
                end
            end
            if (!updated) begin
                sb_addr[sb_size] = addr;
                sb_data[sb_size] = data;
                sb_size          = sb_size + 1;
            end
        end
    endtask

    task automatic sb_check;
        input [24:0] addr;
        input [63:0] data;
        reg          found;
        begin
            found = 1'b0;
            for (sb_idx = 0; sb_idx < sb_size; sb_idx = sb_idx + 1) begin
                if (sb_addr[sb_idx] == addr) begin
                    found = 1'b1;
                    if (sb_data[sb_idx] !== data) begin
                        $display("[%0t] ERROR: addr=%0d expected=0x%016h got=0x%016h",
                                 $time, addr, sb_data[sb_idx], data);
                        $fatal;
                    end
                end
            end
            if (!found) begin
                $display("[%0t] ERROR: read from unknown addr=%0d data=0x%016h",
                         $time, addr, data);
                // Treat reads from never-written locations as fatal in
                // production-style runs so that any unintended access
                // pattern is caught immediately.
                $fatal;
            end
        end
    endtask

    // ------------------------------------------------------------------------
    // Host command sanity: flag illegal CMD encodings at enqueue time and
    // enforce basic FIFO handshake rules (cmd_put only when NOTFULL=1).
    // As in the core-top testbench, the NOTFULL check is tolerant of the
    // single-cycle boundary where FILLCOUNT has just entered the "full" region
    // on the same edge that the host asserts cmd_put based on the previous
    // cycle's NOTFULL=1 observation. Only true overruns (writes beyond the
    // documented safe region) are treated as errors.
    // ------------------------------------------------------------------------
    always @(posedge CLK) begin
        if (cmd_put) begin
            if (CMD !== CMD_NOP &&
                CMD !== CMD_SCR &&
                CMD !== CMD_SCW &&
                CMD !== CMD_BLR &&
                CMD !== CMD_BLW) begin
`ifdef NEGATIVE_TESTS
                if (neg_expect_illegal_cmd) begin
                    // In NEGATIVE_TESTS mode this particular illegal CMD is
                    // expected and treated as a passing condition, so we do
                    // not terminate the simulation here.
                    $display("[%0t] NEG: expected illegal CMD encoding observed: CMD=%0b SZ=%0b ADDR=%0d",
                             $time, CMD, SZ, ADDR);
                end else begin
                    $display("[%0t] ERROR: Host issued illegal CMD encoding: CMD=%0b SZ=%0b ADDR=%0d",
                             $time, CMD, SZ, ADDR);
                    $fatal;
                end
`else
                $display("[%0t] ERROR: Host issued illegal CMD encoding: CMD=%0b SZ=%0b ADDR=%0d",
                         $time, CMD, SZ, ADDR);
                $fatal;
`endif
            end
            if (!NOTFULL && (FILLCOUNT > 7'd33)) begin
                $display("[%0t] ERROR: cmd_put asserted while NOTFULL=0 (host overrun, fillcount=%0d).",
                         $time, FILLCOUNT);
            end
        end
    end

    localparam CLK_PERIOD = 2;   // 500 MHz
    localparam CMD_NOP  = 3'b000;
    localparam CMD_SCR  = 3'b001;
    localparam CMD_SCW  = 3'b010;
    localparam CMD_BLR  = 3'b011;
    localparam CMD_BLW  = 3'b100;

    initial CLK = 0;
    always #(CLK_PERIOD/2) CLK = ~CLK;

    // DUT: server-style wrapper around the core controller.
    ddr2_server_controller u_dut (
        .CLK(CLK),
        .RESET(RESET),
        .INITDDR(INITDDR),
        .CMD(CMD),
        .SZ(SZ),
        .ADDR(ADDR),
        .cmd_put(cmd_put),
        .DIN(DIN),
        .put_dataFIFO(put_dataFIFO),
        .FETCHING(FETCHING),
        .SELFREF_REQ(SELFREF_REQ),
        .SELFREF_EXIT(SELFREF_EXIT),
        .PWRDOWN_REQ(PWRDOWN_REQ),
        .PWRDOWN_EXIT(PWRDOWN_EXIT),
        .DLL_REQ(DLL_REQ),
        .DLL_MODE(DLL_MODE),
        .DOUT(DOUT),
        .RADDR(RADDR),
        .FILLCOUNT(FILLCOUNT),
        .READY(READY),
        .VALIDOUT(VALIDOUT),
        .NOTFULL(NOTFULL),
        .C0_CSBAR_PAD(C0_CSBAR_PAD),
        .C0_RASBAR_PAD(C0_RASBAR_PAD),
        .C0_CASBAR_PAD(C0_CASBAR_PAD),
        .C0_WEBAR_PAD(C0_WEBAR_PAD),
        .C0_BA_PAD(C0_BA_PAD),
        .C0_A_PAD(C0_A_PAD),
        .C0_DM_PAD(C0_DM_PAD),
        .C0_ODT_PAD(C0_ODT_PAD),
        .C0_CK_PAD(C0_CK_PAD),
        .C0_CKBAR_PAD(C0_CKBAR_PAD),
        .C0_CKE_PAD(C0_CKE_PAD),
        .C0_DQ_PAD(C0_DQ_PAD),
        .C0_DQS_PAD(C0_DQS_PAD),
        .C0_DQSBAR_PAD(C0_DQSBAR_PAD)
`ifdef SIM_DIRECT_READ
        ,
        .sim_mem_rd_valid(MEM_RD_VALID),
        .sim_mem_rd_data(MEM_RD_DATA)
`endif
    );

    // Simple behavioral DDR2 memory model connected to the pad interface.
    // Exposes internal read/write activity for closed-loop validation.
    wire        MEM_WR_VALID;
    wire [31:0] MEM_WR_ADDR;
    wire [15:0] MEM_WR_DATA;
    wire        MEM_RD_VALID;
    wire [31:0] MEM_RD_ADDR;
    wire [15:0] MEM_RD_DATA;

    // Allow build-time override of the memory model's parameters (depth, read
    // latency, rank count) so that the same server-top testbench can be reused
    // across multiple logical configurations in regression.
`ifdef MEM_DEPTH_OVERRIDE
    localparam integer MEM_DEPTH_TB  = `MEM_DEPTH_OVERRIDE;
`else
    localparam integer MEM_DEPTH_TB  = 1024;
`endif
`ifdef READ_LAT_OVERRIDE
    localparam integer READ_LAT_TB   = `READ_LAT_OVERRIDE;
`else
    localparam integer READ_LAT_TB   = 24;
`endif
`ifdef RANK_BITS_OVERRIDE
    localparam integer RANK_BITS_TB  = `RANK_BITS_OVERRIDE;
`else
    localparam integer RANK_BITS_TB  = 1;
`endif

    ddr2_simple_mem #(
        .MEM_DEPTH(MEM_DEPTH_TB),
        // Align READ latency with controller's internal SCREAD/SCREND timing
        // so that the model begins driving data while the return path is
        // actively capturing it.
        .READ_LAT(READ_LAT_TB),
        // Two-rank-capable model; its CS# vector is driven directly from the
        // server controller's per-rank CS# outputs.
        .RANK_BITS(RANK_BITS_TB)
    ) u_mem (
        .clk(CLK),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad_vec(C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .ba_pad(C0_BA_PAD),
        .a_pad(C0_A_PAD),
        .dq_pad(C0_DQ_PAD),
        .dqs_pad(C0_DQS_PAD),
        .dqsbar_pad(C0_DQSBAR_PAD),
        .dbg_wr_valid(MEM_WR_VALID),
        .dbg_wr_addr(MEM_WR_ADDR),
        .dbg_wr_data(MEM_WR_DATA),
        .dbg_rd_valid(MEM_RD_VALID),
        .dbg_rd_addr(MEM_RD_ADDR),
        .dbg_rd_data(MEM_RD_DATA)
    );

    // ------------------------------------------------------------------------
    // Protocol / timing monitors (identical to tb_ddr2_controller).
    // ------------------------------------------------------------------------
    ddr2_fifo_monitor u_fifo_mon (
        .clk(CLK),
        .reset(RESET),
        .fillcount(FILLCOUNT),
        .notfull(NOTFULL)
    );

    ddr2_refresh_monitor u_ref_mon (
        .clk(CLK),
        .reset(RESET),
        .ready_i(READY),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD)
    );

    ddr2_timing_checker u_timing_chk (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .ba_pad(C0_BA_PAD)
    );

    // Turnaround / write-or-read-to-precharge timing checker for server top.
    ddr2_turnaround_checker u_turnaround_chk (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad_any(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .ba_pad(C0_BA_PAD)
    );

    ddr2_bank_checker u_bank_chk (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .ba_pad(C0_BA_PAD),
        .a_pad(C0_A_PAD)
    );

    ddr2_dqs_monitor u_dqs_mon (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .dqs_pad(C0_DQS_PAD)
    );

    // OCD / ZQ calibration monitor (server top): same checks as the core-top
    // monitor, connected to the shared DDR2 bus.
    ddr2_ocd_zq_monitor #(
        .EMRS1_OCD_ENTER_VAL(13'h0600),
        .EMRS1_OCD_EXIT_VAL (13'h0640),
        .TOCD_MIN_CYCLES   (10),
        .TZQINIT_MIN_CYCLES(0)
    ) u_ocd_zq_mon (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_pad(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD),
        .ba_pad(C0_BA_PAD),
        .a_pad(C0_A_PAD)
    );

    // Power-mode monitor (server top): mirrors the core-top checker.
    ddr2_power_monitor u_power_mon (
        .clk(CLK),
        .reset(RESET),
        .cke_pad(C0_CKE_PAD),
        .csbar_any(&C0_CSBAR_PAD),
        .rasbar_pad(C0_RASBAR_PAD),
        .casbar_pad(C0_CASBAR_PAD),
        .webar_pad(C0_WEBAR_PAD)
    );

`ifndef SIM_DIRECT_READ
    // Closed-loop checks (full bus-level mode), as in tb_ddr2_controller.
    reg [15:0] last_mem_rd_data;
    reg        mem_rd_seen;

    always @(posedge CLK) begin
        if (RESET) begin
            last_mem_rd_data <= 16'h0000;
            mem_rd_seen      <= 1'b0;
        end else begin
            if (MEM_RD_VALID) begin
                last_mem_rd_data <= MEM_RD_DATA;
                mem_rd_seen      <= 1'b1;
            end
            if (VALIDOUT && !mem_rd_seen) begin
                $display("[%0t] ERROR: VALIDOUT asserted before any MEM_RD_VALID.",
                         $time);
                $fatal;
            end
        end
    end
`endif

    // ------------------------------------------------------------------------
    // Helper tasks (mostly identical to tb_ddr2_controller).
    // ------------------------------------------------------------------------
    task automatic do_scalar_rw;
        input [24:0] addr;
        reg   [15:0] data16;
        reg   [63:0] data64;
        begin
            data16 = pattern_for_addr(addr);
            // Replicate the 16-bit pattern across all four lanes so that each
            // slice sees identical data for this address.
            data64 = {4{data16}};

            @(posedge CLK);
            while (!NOTFULL) begin
                @(posedge CLK);
            end
            ADDR         = addr;
            CMD          = CMD_SCW;
            SZ           = 2'b00;
            cmd_put      = 1'b1;
            DIN          = data64;
            put_dataFIFO = 1'b1;
            @(posedge CLK);
            cmd_put      = 1'b0;
            put_dataFIFO = 1'b0;
            $display("[%0t] SCW issued (server): addr=%0d data16=0x%04h", $time, addr, data16);

            sb_write(addr, data64);

            repeat (200) @(posedge CLK);

            @(posedge CLK);
            CMD     = CMD_SCR;
            SZ      = 2'b00;
            ADDR    = addr;
            cmd_put = 1'b1;
            @(posedge CLK);
            cmd_put = 1'b0;
            $display("[%0t] SCR issued: addr=%0d", $time, addr);

            FETCHING = 1'b1;
            wait (VALIDOUT === 1'b1);
            @(posedge CLK);

            FETCHING = 1'b0;
            repeat (50) @(posedge CLK);
        end
    endtask

    task automatic do_block_rw;
        input [24:0] base_addr;
        input [1:0]  sz;
        integer      nwords;
        integer      beat;
        integer      wait_cycles;
        reg [15:0]  data16;
        reg [63:0]  data64;
        begin
            case (sz)
                2'b00: nwords = 8;
                2'b01: nwords = 16;
                2'b10: nwords = 24;
                2'b11: nwords = 32;
                default: nwords = 8;
            endcase

            @(posedge CLK);
            while (!NOTFULL) begin
                @(posedge CLK);
            end

            ADDR    = base_addr;
            CMD     = CMD_BLW;
            SZ      = sz;
            cmd_put = 1'b1;
            @(posedge CLK);
            cmd_put = 1'b0;
            $display("[%0t] BLW issued: base_addr=%0d SZ=%0d (nwords=%0d)",
                     $time, base_addr, sz, nwords);

            for (beat = 0; beat < nwords; beat = beat + 1) begin
                data16       = pattern_for_addr(base_addr + beat[24:0]);
                data64       = {4{data16}};
                DIN          = data64;
                put_dataFIFO = 1'b1;
                @(posedge CLK);
                put_dataFIFO = 1'b0;
                @(posedge CLK);
                sb_write(base_addr + beat[24:0], data64);
            end

            repeat (600) @(posedge CLK);

            @(posedge CLK);
            ADDR    = base_addr;
            CMD     = CMD_BLR;
            SZ      = sz;
            cmd_put = 1'b1;
            @(posedge CLK);
            cmd_put = 1'b0;
            $display("[%0t] BLR issued: base_addr=%0d SZ=%0d (expect %0d beats)",
                     $time, base_addr, sz, nwords);

            FETCHING    = 1'b1;
            beat        = 0;
            wait_cycles = 0;
`ifdef SIM_DIRECT_READ
            while (beat < nwords) begin
                @(posedge CLK);
                wait_cycles = wait_cycles + 1;
                if (VALIDOUT) begin
                    $display("[%0t] BLR beat %0d observed: RADDR=%0d DOUT=0x%04h",
                             $time, beat, RADDR, DOUT);
                    beat        = beat + 1;
                    wait_cycles = 0;
                end
                if (wait_cycles > 20000) begin
                    $display("[%0t] FATAL: BLR timeout waiting for beat %0d/%0d (VALIDOUT stuck low).",
                             $time, beat, nwords);
                    $fatal;
                end
            end
`else
            while (wait_cycles <= 20000) begin
                @(posedge CLK);
                wait_cycles = wait_cycles + 1;
                if (VALIDOUT) begin
                    $display("[%0t] BLR beat (bus mode) observed: RADDR=%0d DOUT=0x%04h",
                             $time, RADDR, DOUT);
                    wait_cycles = 0;
                end
            end
`endif

            $display("[%0t] BLW/BLR sequence OK: base_addr=%0d SZ=%0d (nwords=%0d)",
                     $time, base_addr, sz, nwords);

            FETCHING = 1'b0;
            repeat (100) @(posedge CLK);
        end
    endtask

    // Ranked variants: encode a logical rank into the MSB of ADDR so that the
    // server controller's internal RANK_SEL hint and two-rank CS# steering are
    // exercised while reusing the existing helper behavior.
    task automatic do_scalar_rw_ranked;
        input [24:0] addr;
        input        rank;
        reg   [24:0] addr_full;
        begin
            addr_full = {rank, addr[23:0]};
            do_scalar_rw(addr_full);
        end
    endtask

    task automatic do_block_rw_ranked;
        input [24:0] base_addr;
        input [1:0]  sz;
        input        rank;
        reg   [24:0] base_full;
        begin
            base_full = {rank, base_addr[23:0]};
            do_block_rw(base_full, sz);
        end
    endtask

    task automatic do_scalar_read_uninitialized;
        input [24:0] addr;
        begin
            @(posedge CLK);
            while (!NOTFULL) begin
                @(posedge CLK);
            end
            ADDR    = addr;
            CMD     = CMD_SCR;
            SZ      = 2'b00;
            cmd_put = 1'b1;
            @(posedge CLK);
            cmd_put = 1'b0;
            $display("[%0t] NEG: SCR (no prior write) issued: addr=%0d", $time, addr);

            FETCHING = 1'b1;
            wait (VALIDOUT === 1'b1);
            @(posedge CLK);
            FETCHING = 1'b0;
        end
    endtask

    task automatic run_random_traffic;
        integer n_iter;
        integer choice;
        reg [24:0] rand_addr;
        reg [1:0]  rand_sz;
        begin
            $display("[%0t] Starting randomized traffic phase (server top)...", $time);
            rand_addr = 25'd0;

            for (n_iter = 0; n_iter < 64; n_iter = n_iter + 1) begin
                /* verilator lint_off WIDTHTRUNC */
                rand_addr = $urandom % 1024;
                rand_sz   = $urandom % 4;
                /* verilator lint_on WIDTHTRUNC */
                choice    = $urandom % 4;
                case (choice)
                    0: do_scalar_rw(rand_addr);
                    1: do_block_rw(rand_addr & 25'hFFFFF8, 2'b00);
                    default: do_block_rw(rand_addr & 25'hFFFFF8, rand_sz);
                endcase
            end

            $display("[%0t] Randomized traffic phase (server top) completed.", $time);
        end
    endtask

    // ------------------------------------------------------------------------
    // Monitor / main stimulus (mostly identical to tb_ddr2_controller).
    // ------------------------------------------------------------------------
    always @(posedge CLK) begin
`ifdef CSV_TRACE
        $fwrite(csv_fd,
                "%0t,%0d,%0d,%0d,%0d,%0b,%0b,%0h,%0d,%0b,%0d,%0h,%0b,%0d,%0h\n",
                $time, cycle,
                CMD, SZ, ADDR,
                FETCHING, VALIDOUT, DOUT, RADDR,
                MEM_WR_VALID, MEM_WR_ADDR, MEM_WR_DATA,
                MEM_RD_VALID, MEM_RD_ADDR, MEM_RD_DATA);
`endif

        if (!C0_CSBAR_PAD && !C0_RASBAR_PAD && !C0_CASBAR_PAD && C0_WEBAR_PAD) begin
            $display("[%0t] Detected AUTO REFRESH command on DDR2 bus (server top).", $time);
        end

        if (cmd_put) begin
            case (CMD)
                CMD_SCW: cov_scw <= cov_scw + 1;
                CMD_SCR: cov_scr <= cov_scr + 1;
                CMD_BLW: cov_blw <= cov_blw + 1;
                CMD_BLR: cov_blr <= cov_blr + 1;
                default: ;
            endcase
            case (SZ)
                2'b00: cov_sz0 <= cov_sz0 + 1;
                2'b01: cov_sz1 <= cov_sz1 + 1;
                2'b10: cov_sz2 <= cov_sz2 + 1;
                2'b11: cov_sz3 <= cov_sz3 + 1;
            endcase
        end

        if (VALIDOUT) begin
            $display("[%0t] READ observed (server top): RADDR=%0d DOUT=0x%016h", $time, RADDR, DOUT);
`ifdef SIM_DIRECT_READ
            sb_check(RADDR, DOUT);
`endif
        end
    end

    initial begin
        $dumpfile("tb_ddr2_server_controller.iverilog.vcd");
        $dumpvars(0, tb_ddr2_server_controller);
        cycle = 0;
`ifdef NEGATIVE_TESTS
        neg_expect_illegal_cmd = 1'b0;
`endif
`ifdef CSV_TRACE
        csv_fd = $fopen("ddr2_trace_server.csv", "w");
        $fwrite(csv_fd, "time,cycle,CMD,SZ,ADDR,FETCHING,VALIDOUT,DOUT,RADDR,MEM_WR_VALID,MEM_WR_ADDR,MEM_WR_DATA,MEM_RD_VALID,MEM_RD_ADDR,MEM_RD_DATA\n");
`endif
        RESET    = 1;
        INITDDR  = 0;
        CMD      = CMD_NOP;
        SZ       = 2'b00;
        ADDR     = 25'b0;
        cmd_put  = 0;
        DIN      = 64'b0;
        put_dataFIFO = 0;
        FETCHING = 0;
        SELFREF_REQ  = 0;
        SELFREF_EXIT = 0;
        PWRDOWN_REQ  = 0;
        PWRDOWN_EXIT = 0;
        DLL_REQ      = 0;
        DLL_MODE     = 0;
        SELFREF_REQ  = 0;
        SELFREF_EXIT = 0;
        PWRDOWN_REQ  = 0;
        PWRDOWN_EXIT = 0;
        repeat (10) @(posedge CLK);
        RESET = 0;
        @(posedge CLK);
        INITDDR = 1;
        @(posedge CLK);
        INITDDR = 0;
        $display("[%0t] (server) INITDDR asserted, waiting for READY...", $time);
        while (!READY) begin
            @(posedge CLK);
            cycle = cycle + 1;
            if (cycle % 20000 == 0 && cycle > 0)
                $display("[%0t] (server) cycle %0d, READY=%b", $time, cycle, READY);
        end
        $display("[%0t] (server) READY asserted at cycle %0d", $time, cycle);

        @(posedge CLK);
        if (NOTFULL)
            $display("[%0t] (server) NOTFULL=1 (FIFOs can accept commands)", $time);
        else
            $display("[%0t] (server) NOTFULL=0", $time);

        sb_reset();

        cov_scw = 0;
        cov_scr = 0;
        cov_blw = 0;
        cov_blr = 0;
        cov_sz0 = 0;
        cov_sz1 = 0;
        cov_sz2 = 0;
        cov_sz3 = 0;

        // Reuse the same scenario set as tb_ddr2_controller.
        do_scalar_rw(25'd0);
        do_scalar_rw(25'd1);
        do_scalar_rw(25'd128);
        do_scalar_rw(25'd512);

        do_block_rw(25'd32,   2'b00);
        do_block_rw(25'd256,  2'b01);
        do_block_rw(25'd384,  2'b10);
        do_block_rw(25'd512,  2'b11);

        $display("[%0t] (server) Starting FIFO stress / refresh-interleaving test...", $time);
        for (i = 0; i < 8; i = i + 1) begin
            do_scalar_rw(25'd600 + i[24:0]);
            /* verilator lint_off WIDTHTRUNC */
            do_block_rw(700 + (i * 40), 2'b01);
            /* verilator lint_on WIDTHTRUNC */
        end

        $display("[%0t] (server) Starting reset-during-traffic robustness test...", $time);
        do_scalar_rw(25'd900);
        do_block_rw(25'd920, 2'b00);

        $display("[%0t] (server) Asserting RESET in the middle of activity...", $time);
        RESET    = 1'b1;
        INITDDR  = 1'b0;
        CMD      = CMD_NOP;
        SZ       = 2'b00;
        ADDR     = 25'b0;
        cmd_put  = 1'b0;
        DIN      = 64'b0;
        put_dataFIFO = 1'b0;
        FETCHING = 1'b0;
        repeat (10) @(posedge CLK);

        RESET   = 1'b0;
        @(posedge CLK);
        INITDDR = 1'b1;
        @(posedge CLK);
        INITDDR = 1'b0;
        $display("[%0t] (server) Re-INITDDR asserted after mid-traffic reset, waiting for READY...", $time);
        cycle = 0;
        while (!READY) begin
            @(posedge CLK);
            cycle = cycle + 1;
            if (cycle % 20000 == 0 && cycle > 0)
                $display("[%0t] (server post-reset) cycle %0d, READY=%b", $time, cycle, READY);
        end
        $display("[%0t] (server) READY re-asserted after reset at cycle %0d", $time, cycle);

        sb_reset();
        do_scalar_rw(25'd32);
        do_block_rw(25'd64, 2'b01);

        // --------------------------------------------------------------------
        // Manual self-refresh and precharge power-down (server top)
        // --------------------------------------------------------------------
        $display("[%0t] (server) Starting manual self-refresh / power-down tests...", $time);

        // Ensure the front-end is idle before requesting self-refresh.
        @(posedge CLK);
        while (!READY || !NOTFULL) begin
            @(posedge CLK);
        end

        $display("[%0t] (server) Asserting SELFREF_REQ...", $time);
        SELFREF_REQ = 1'b1;
        @(posedge CLK);
        SELFREF_REQ = 1'b0;

        // Hold self-refresh for a while.
        repeat (2000) @(posedge CLK);

        $display("[%0t] (server) Asserting SELFREF_EXIT...", $time);
        SELFREF_EXIT = 1'b1;
        @(posedge CLK);
        SELFREF_EXIT = 1'b0;
        repeat (2000) @(posedge CLK);

        // Sanity-check: scalar/block traffic after exit.
        sb_reset();
        do_scalar_rw(25'd40);
        do_block_rw(25'd72, 2'b00);

        // Precharge power-down sequence.
        @(posedge CLK);
        while (!READY || !NOTFULL) begin
            @(posedge CLK);
        end

        $display("[%0t] (server) Asserting PWRDOWN_REQ...", $time);
        PWRDOWN_REQ = 1'b1;
        @(posedge CLK);
        PWRDOWN_REQ = 1'b0;

        repeat (2000) @(posedge CLK);

        $display("[%0t] (server) Asserting PWRDOWN_EXIT...", $time);
        PWRDOWN_EXIT = 1'b1;
        @(posedge CLK);
        PWRDOWN_EXIT = 1'b0;
        repeat (1000) @(posedge CLK);

        sb_reset();
        do_scalar_rw(25'd96);
        do_block_rw(25'd128, 2'b01);

        // --------------------------------------------------------------------
        // Multi-rank bus-level exercise (server top)
        // - Encode a logical rank into the MSB of ADDR so that the server
        //   wrapper's RANK_SEL hint and two-rank CS# steering are both
        //   exercised through the shared DDR2 bus and memory model.
        // --------------------------------------------------------------------
        $display("[%0t] (server) Starting multi-rank bus-level exercise (rank 0 vs rank 1)...", $time);
        // Scalar traffic to the same low addresses but different rank bits.
        do_scalar_rw_ranked(25'd32,  1'b0);
        do_scalar_rw_ranked(25'd32,  1'b1);
        do_scalar_rw_ranked(25'd128, 1'b0);
        do_scalar_rw_ranked(25'd128, 1'b1);

        // Block traffic to identical base addresses on two logical ranks.
        do_block_rw_ranked(25'd256, 2'b00, 1'b0);
        do_block_rw_ranked(25'd256, 2'b00, 1'b1);

        run_random_traffic();

        repeat (2000) @(posedge CLK);

        $display("----------------------------------------------------------------");
        $display("DDR2 SERVER controller functional coverage (approximate):");
        $display("  SCW count = %0d", cov_scw);
        $display("  SCR count = %0d", cov_scr);
        $display("  BLW count = %0d", cov_blw);
        $display("  BLR count = %0d", cov_blr);
        $display("  SZ=00 count = %0d", cov_sz0);
        $display("  SZ=01 count = %0d", cov_sz1);
        $display("  SZ=10 count = %0d", cov_sz2);
        $display("  SZ=11 count = %0d", cov_sz3);
        $display("----------------------------------------------------------------");

        $display("[%0t] (server) All tests completed successfully.", $time);

`ifdef NEGATIVE_TESTS
        $display("[%0t] (server) Starting NEGATIVE_TESTS...", $time);
        @(posedge CLK);
        while (!NOTFULL) begin
            @(posedge CLK);
        end
        neg_expect_illegal_cmd = 1'b1;
        ADDR    = 25'd16;
        CMD     = 3'b111;
        SZ      = 2'b00;
        cmd_put = 1'b1;
        @(posedge CLK);
        cmd_put = 1'b0;
        neg_expect_illegal_cmd = 1'b0;
        $display("[%0t] (server) NEG: illegal CMD=3'b111 enqueued.", $time);
        // do_scalar_read_uninitialized(25'd1023);
`endif
`ifdef CSV_TRACE
        $fclose(csv_fd);
`endif
        $finish;
    end

endmodule
/* verilator lint_on UNUSEDSIGNAL */

